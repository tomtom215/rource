(* SPDX-License-Identifier: GPL-3.0-or-later *)
(* Copyright (C) 2026 Tom F <https://github.com/tomtom215> *)

(**
 * RourceMath_Extract.v - Unified Coq Extraction for All rource-math Types
 *
 * This module extracts ALL computational types (ZVec2, ZVec3, ZVec4,
 * ZMat3, ZMat4, ZColor, ZRect, zlerp, zclamp) into a single OCaml
 * module. This unified extraction
 * is the input for the Coq-to-WASM pipeline:
 *
 *   RourceMath_Extract.v (this file)
 *     │
 *     ▼  [Coq Standard Extraction]
 *   rource_math_extracted.ml (OCaml)
 *     │
 *     ▼  [ocamlfind ocamlc / wasm_of_ocaml]
 *   rource_math.wasm (WebAssembly)
 *
 * VERIFICATION STATUS: PEER REVIEWED PUBLISHED ACADEMIC STANDARD
 * - All source types have zero admits
 * - Combined: 8 types, 160+ theorems proven across all Compute files
 * - Extraction is semantics-preserving (Coq guarantee)
 *)

Require Import ZArith.
Require Import ExtrOcamlBasic.
Require Import ExtrOcamlZInt.

Set Warnings "-notation-overridden".
Require Import RourceMath.Vec2_Compute.
Require Import RourceMath.Vec3_Compute.
Require Import RourceMath.Vec4_Compute.
Require Import RourceMath.Mat3_Compute.
Require Import RourceMath.Mat4_Compute.
Require Import RourceMath.Color_Compute.
Require Import RourceMath.Rect_Compute.
Require Import RourceMath.Utils_Compute.
Set Warnings "default".

(** * Unified Extraction *)

Extraction "rource_math_extracted"
  (* Vec2 *)
  ZVec2 mkZVec2 zvec2_x zvec2_y
  zvec2_new zvec2_zero zvec2_splat zvec2_unit_x zvec2_unit_y
  zvec2_add zvec2_sub zvec2_neg zvec2_scale zvec2_mul
  zvec2_dot zvec2_cross zvec2_perp zvec2_length_squared
  zvec2_eq_dec
  (* Vec3 *)
  ZVec3 mkZVec3 zvec3_x zvec3_y zvec3_z
  zvec3_new zvec3_zero zvec3_splat zvec3_unit_x zvec3_unit_y zvec3_unit_z
  zvec3_add zvec3_sub zvec3_neg zvec3_scale zvec3_mul
  zvec3_dot zvec3_cross zvec3_length_squared zvec3_scalar_triple
  zvec3_eq_dec
  (* Vec4 *)
  ZVec4 mkZVec4 zvec4_x zvec4_y zvec4_z zvec4_w
  zvec4_new zvec4_zero zvec4_one zvec4_splat
  zvec4_unit_x zvec4_unit_y zvec4_unit_z zvec4_unit_w
  zvec4_add zvec4_sub zvec4_neg zvec4_scale zvec4_mul
  zvec4_dot zvec4_length_squared
  zvec4_eq_dec
  (* Mat3 *)
  ZMat3 mkZMat3 zm3_0 zm3_1 zm3_2 zm3_3 zm3_4 zm3_5 zm3_6 zm3_7 zm3_8
  zmat3_zero zmat3_identity zmat3_add zmat3_neg zmat3_sub
  zmat3_scale zmat3_transpose zmat3_mul zmat3_determinant zmat3_trace
  (* Mat4 *)
  ZMat4 mkZMat4
  zm4_0 zm4_1 zm4_2 zm4_3 zm4_4 zm4_5 zm4_6 zm4_7
  zm4_8 zm4_9 zm4_10 zm4_11 zm4_12 zm4_13 zm4_14 zm4_15
  zmat4_zero zmat4_identity zmat4_add zmat4_neg zmat4_sub
  zmat4_scale zmat4_transpose zmat4_mul zmat4_trace
  (* Color *)
  ZColor mkZColor zcolor_r zcolor_g zcolor_b zcolor_a
  zcolor_new zcolor_rgb zcolor_gray zcolor_transparent zcolor_black zcolor_white
  zcolor_with_alpha zcolor_fade zcolor_lerp zcolor_premultiplied
  zcolor_blend_over zcolor_luminance zcolor_clamp zcolor_eq_dec
  (* Rect *)
  ZRect mkZRect zrect_x zrect_y zrect_w zrect_h
  zrect_new zrect_zero zrect_right zrect_bottom zrect_area zrect_perimeter
  zrect_center_x zrect_center_y zrect_is_valid zrect_is_empty
  zrect_contains_point zrect_contains_rect zrect_intersects
  zrect_translate zrect_expand zrect_shrink zrect_union zrect_eq_dec
  (* Utils *)
  zlerp zclamp.
