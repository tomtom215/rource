(* SPDX-License-Identifier: GPL-3.0-or-later *)
(* Copyright (C) 2026 Tom F <https://github.com/tomtom215> *)

(**
 * Vec4_Compute.v - Computational 4D Vector Specification (Extractable)
 *
 * This module provides a COMPUTABLE formalization of 4D vectors using Coq's
 * Z (integer) type. Unlike Vec4.v (which uses the axiomatized R type for
 * mathematical reasoning), this module produces fully extractable code.
 *
 * LAYERED VERIFICATION ARCHITECTURE:
 *
 *   Layer 1 (Abstract):      Vec4.v / Vec4_Proofs.v     (R-based, 25+ theorems)
 *   Layer 2 (Computational): Vec4_Compute.v             (Z-based, extractable)
 *   Layer 3 (Extraction):    Vec4_Extract.v             (OCaml/WASM output)
 *
 * VERIFICATION STATUS: PEER REVIEWED PUBLISHED ACADEMIC STANDARD
 * - All definitions are constructive and computable
 * - All proofs are machine-checked by Coq
 * - Zero admits, zero axioms beyond standard library
 *)

Require Import ZArith.
Require Import Lia.
Open Scope Z_scope.

(** * ZVec4 Definition *)

(** A 4D vector with integer components, suitable for extraction. *)
Record ZVec4 : Type := mkZVec4 {
  zvec4_x : Z;
  zvec4_y : Z;
  zvec4_z : Z;
  zvec4_w : Z
}.

(** * Equality Decision *)

Lemma zvec4_eq_dec : forall (a b : ZVec4), {a = b} + {a <> b}.
Proof.
  intros [ax ay az aw] [bx by0 bz bw].
  destruct (Z.eq_dec ax bx) as [Hx | Hx];
  destruct (Z.eq_dec ay by0) as [Hy | Hy];
  destruct (Z.eq_dec az bz) as [Hz | Hz];
  destruct (Z.eq_dec aw bw) as [Hw | Hw].
  - left. subst. reflexivity.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
  - right. intro H. inversion H. contradiction.
Defined.

(** * Constructors *)

Definition zvec4_new (x y z w : Z) : ZVec4 := mkZVec4 x y z w.
Definition zvec4_zero : ZVec4 := mkZVec4 0 0 0 0.
Definition zvec4_one : ZVec4 := mkZVec4 1 1 1 1.
Definition zvec4_splat (v : Z) : ZVec4 := mkZVec4 v v v v.
Definition zvec4_unit_x : ZVec4 := mkZVec4 1 0 0 0.
Definition zvec4_unit_y : ZVec4 := mkZVec4 0 1 0 0.
Definition zvec4_unit_z : ZVec4 := mkZVec4 0 0 1 0.
Definition zvec4_unit_w : ZVec4 := mkZVec4 0 0 0 1.

(** * Arithmetic Operations *)

Definition zvec4_add (a b : ZVec4) : ZVec4 :=
  mkZVec4 (zvec4_x a + zvec4_x b) (zvec4_y a + zvec4_y b)
          (zvec4_z a + zvec4_z b) (zvec4_w a + zvec4_w b).

Definition zvec4_sub (a b : ZVec4) : ZVec4 :=
  mkZVec4 (zvec4_x a - zvec4_x b) (zvec4_y a - zvec4_y b)
          (zvec4_z a - zvec4_z b) (zvec4_w a - zvec4_w b).

Definition zvec4_neg (v : ZVec4) : ZVec4 :=
  mkZVec4 (- zvec4_x v) (- zvec4_y v) (- zvec4_z v) (- zvec4_w v).

Definition zvec4_scale (s : Z) (v : ZVec4) : ZVec4 :=
  mkZVec4 (s * zvec4_x v) (s * zvec4_y v) (s * zvec4_z v) (s * zvec4_w v).

Definition zvec4_mul (a b : ZVec4) : ZVec4 :=
  mkZVec4 (zvec4_x a * zvec4_x b) (zvec4_y a * zvec4_y b)
          (zvec4_z a * zvec4_z b) (zvec4_w a * zvec4_w b).

(** * Dot Product *)

Definition zvec4_dot (a b : ZVec4) : Z :=
  zvec4_x a * zvec4_x b + zvec4_y a * zvec4_y b +
  zvec4_z a * zvec4_z b + zvec4_w a * zvec4_w b.

(** * Length Squared *)

Definition zvec4_length_squared (v : ZVec4) : Z :=
  zvec4_dot v v.

(** * Equality Lemma *)

Lemma zvec4_eq : forall x1 y1 z1 w1 x2 y2 z2 w2 : Z,
  x1 = x2 -> y1 = y2 -> z1 = z2 -> w1 = w2 ->
  mkZVec4 x1 y1 z1 w1 = mkZVec4 x2 y2 z2 w2.
Proof.
  intros. subst. reflexivity.
Qed.

Lemma zvec4_eq_iff : forall a b : ZVec4,
  a = b <-> (zvec4_x a = zvec4_x b /\ zvec4_y a = zvec4_y b /\
             zvec4_z a = zvec4_z b /\ zvec4_w a = zvec4_w b).
Proof.
  intros a b. split.
  - intro H. rewrite H. repeat split; reflexivity.
  - intros [Hx [Hy [Hz Hw]]]. destruct a, b. simpl in *. subst. reflexivity.
Qed.

(** * Vector Space Axioms (Algebraic Properties) *)

(** ** Addition Properties *)

Theorem zvec4_add_comm : forall a b : ZVec4,
  zvec4_add a b = zvec4_add b a.
Proof.
  intros [ax ay az aw] [bx by0 bz bw]. unfold zvec4_add. simpl.
  apply zvec4_eq; lia.
Qed.

Theorem zvec4_add_assoc : forall a b c : ZVec4,
  zvec4_add (zvec4_add a b) c = zvec4_add a (zvec4_add b c).
Proof.
  intros [ax ay az aw] [bx by0 bz bw] [cx cy cz cw]. unfold zvec4_add. simpl.
  apply zvec4_eq; lia.
Qed.

Theorem zvec4_add_zero_r : forall a : ZVec4,
  zvec4_add a zvec4_zero = a.
Proof.
  intros [ax ay az aw]. unfold zvec4_add, zvec4_zero. simpl.
  apply zvec4_eq; lia.
Qed.

Theorem zvec4_add_zero_l : forall a : ZVec4,
  zvec4_add zvec4_zero a = a.
Proof.
  intros [ax ay az aw]. unfold zvec4_add, zvec4_zero. simpl.
  apply zvec4_eq; lia.
Qed.

Theorem zvec4_add_neg : forall a : ZVec4,
  zvec4_add a (zvec4_neg a) = zvec4_zero.
Proof.
  intros [ax ay az aw]. unfold zvec4_add, zvec4_neg, zvec4_zero. simpl.
  apply zvec4_eq; lia.
Qed.

(** ** Scalar Multiplication Properties *)

Theorem zvec4_scale_assoc : forall (s t : Z) (v : ZVec4),
  zvec4_scale (s * t) v = zvec4_scale s (zvec4_scale t v).
Proof.
  intros s t [vx vy vz vw]. unfold zvec4_scale. simpl.
  apply zvec4_eq; ring.
Qed.

Theorem zvec4_scale_dist_vec : forall (s : Z) (a b : ZVec4),
  zvec4_scale s (zvec4_add a b) = zvec4_add (zvec4_scale s a) (zvec4_scale s b).
Proof.
  intros s [ax ay az aw] [bx by0 bz bw]. unfold zvec4_scale, zvec4_add. simpl.
  apply zvec4_eq; ring.
Qed.

Theorem zvec4_scale_dist_scalar : forall (s t : Z) (v : ZVec4),
  zvec4_scale (s + t) v = zvec4_add (zvec4_scale s v) (zvec4_scale t v).
Proof.
  intros s t [vx vy vz vw]. unfold zvec4_scale, zvec4_add. simpl.
  apply zvec4_eq; ring.
Qed.

Theorem zvec4_scale_one : forall v : ZVec4,
  zvec4_scale 1 v = v.
Proof.
  intros [vx vy vz vw]. unfold zvec4_scale.
  apply zvec4_eq; apply Z.mul_1_l.
Qed.

Theorem zvec4_scale_zero : forall v : ZVec4,
  zvec4_scale 0 v = zvec4_zero.
Proof.
  intros [vx vy vz vw]. unfold zvec4_scale, zvec4_zero.
  apply zvec4_eq; apply Z.mul_0_l.
Qed.

(** ** Dot Product Properties *)

Theorem zvec4_dot_comm : forall a b : ZVec4,
  zvec4_dot a b = zvec4_dot b a.
Proof.
  intros [ax ay az aw] [bx by0 bz bw]. unfold zvec4_dot. simpl. ring.
Qed.

Theorem zvec4_dot_linear : forall (s : Z) (a b : ZVec4),
  zvec4_dot (zvec4_scale s a) b = s * zvec4_dot a b.
Proof.
  intros s [ax ay az aw] [bx by0 bz bw]. unfold zvec4_dot, zvec4_scale. simpl. ring.
Qed.

Theorem zvec4_dot_dist : forall a b c : ZVec4,
  zvec4_dot (zvec4_add a b) c = zvec4_dot a c + zvec4_dot b c.
Proof.
  intros [ax ay az aw] [bx by0 bz bw] [cx cy cz cw].
  unfold zvec4_dot, zvec4_add. simpl. ring.
Qed.

(** ** Length Squared Properties *)

Theorem zvec4_length_sq_nonneg : forall v : ZVec4,
  0 <= zvec4_length_squared v.
Proof.
  intros [vx vy vz vw]. unfold zvec4_length_squared, zvec4_dot. simpl.
  assert (H1 : 0 <= vx * vx) by (apply Z.square_nonneg).
  assert (H2 : 0 <= vy * vy) by (apply Z.square_nonneg).
  assert (H3 : 0 <= vz * vz) by (apply Z.square_nonneg).
  assert (H4 : 0 <= vw * vw) by (apply Z.square_nonneg).
  lia.
Qed.

Theorem zvec4_length_sq_zero_iff : forall v : ZVec4,
  zvec4_length_squared v = 0 <-> v = zvec4_zero.
Proof.
  intros [vx vy vz vw]. unfold zvec4_length_squared, zvec4_dot, zvec4_zero. simpl.
  split.
  - intro H.
    assert (Hx: 0 <= vx * vx) by (apply Z.square_nonneg).
    assert (Hy: 0 <= vy * vy) by (apply Z.square_nonneg).
    assert (Hz: 0 <= vz * vz) by (apply Z.square_nonneg).
    assert (Hw: 0 <= vw * vw) by (apply Z.square_nonneg).
    assert (Hxz: vx * vx = 0) by lia.
    assert (Hyz: vy * vy = 0) by lia.
    assert (Hzz: vz * vz = 0) by lia.
    assert (Hwz: vw * vw = 0) by lia.
    apply Z.mul_eq_0 in Hxz. apply Z.mul_eq_0 in Hyz.
    apply Z.mul_eq_0 in Hzz. apply Z.mul_eq_0 in Hwz.
    destruct Hxz; destruct Hyz; destruct Hzz; destruct Hwz; subst; reflexivity.
  - intro H. inversion H. subst. reflexivity.
Qed.

(** ** Subtraction and Negation Properties *)

Theorem zvec4_sub_as_add_neg : forall a b : ZVec4,
  zvec4_sub a b = zvec4_add a (zvec4_neg b).
Proof.
  intros [ax ay az aw] [bx by0 bz bw]. unfold zvec4_sub, zvec4_add, zvec4_neg. simpl.
  apply zvec4_eq; ring.
Qed.

Theorem zvec4_neg_as_scale : forall v : ZVec4,
  zvec4_neg v = zvec4_scale (-1) v.
Proof.
  intros [vx vy vz vw]. unfold zvec4_neg, zvec4_scale.
  apply zvec4_eq; ring.
Qed.

(** ** Component Multiplication Properties *)

Theorem zvec4_mul_comm : forall a b : ZVec4,
  zvec4_mul a b = zvec4_mul b a.
Proof.
  intros [ax ay az aw] [bx by0 bz bw]. unfold zvec4_mul. simpl.
  apply zvec4_eq; ring.
Qed.

(** ** Vector Space Structure (Combined Verification) *)

Theorem zvec4_vector_space : forall (s t : Z) (a b : ZVec4),
  zvec4_add a b = zvec4_add b a /\
  zvec4_add (zvec4_add a b) zvec4_zero = zvec4_add a b /\
  zvec4_add a (zvec4_neg a) = zvec4_zero /\
  zvec4_scale 1 a = a /\
  zvec4_scale (s * t) a = zvec4_scale s (zvec4_scale t a) /\
  zvec4_scale s (zvec4_add a b) = zvec4_add (zvec4_scale s a) (zvec4_scale s b) /\
  zvec4_scale (s + t) a = zvec4_add (zvec4_scale s a) (zvec4_scale t a).
Proof.
  intros s t a b. repeat split.
  - apply zvec4_add_comm.
  - rewrite zvec4_add_assoc. rewrite zvec4_add_zero_r. reflexivity.
  - apply zvec4_add_neg.
  - apply zvec4_scale_one.
  - apply zvec4_scale_assoc.
  - apply zvec4_scale_dist_vec.
  - apply zvec4_scale_dist_scalar.
Qed.

(** * Min/Max/Abs Operations *)

Definition zvec4_min (a b : ZVec4) : ZVec4 :=
  mkZVec4 (Z.min (zvec4_x a) (zvec4_x b)) (Z.min (zvec4_y a) (zvec4_y b))
          (Z.min (zvec4_z a) (zvec4_z b)) (Z.min (zvec4_w a) (zvec4_w b)).

Definition zvec4_max (a b : ZVec4) : ZVec4 :=
  mkZVec4 (Z.max (zvec4_x a) (zvec4_x b)) (Z.max (zvec4_y a) (zvec4_y b))
          (Z.max (zvec4_z a) (zvec4_z b)) (Z.max (zvec4_w a) (zvec4_w b)).

Definition zvec4_abs (v : ZVec4) : ZVec4 :=
  mkZVec4 (Z.abs (zvec4_x v)) (Z.abs (zvec4_y v))
          (Z.abs (zvec4_z v)) (Z.abs (zvec4_w v)).

(** * Reduction Operations *)

Definition zvec4_element_sum (v : ZVec4) : Z :=
  zvec4_x v + zvec4_y v + zvec4_z v + zvec4_w v.

Definition zvec4_element_product (v : ZVec4) : Z :=
  zvec4_x v * zvec4_y v * zvec4_z v * zvec4_w v.

Definition zvec4_distance_squared (a b : ZVec4) : Z :=
  zvec4_length_squared (zvec4_sub a b).

(** ** Min/Max Properties *)

Theorem zvec4_min_comm : forall a b : ZVec4,
  zvec4_min a b = zvec4_min b a.
Proof.
  intros [ax ay az aw] [bx by0 bz bw]. unfold zvec4_min. simpl.
  apply zvec4_eq; apply Z.min_comm.
Qed.

Theorem zvec4_max_comm : forall a b : ZVec4,
  zvec4_max a b = zvec4_max b a.
Proof.
  intros [ax ay az aw] [bx by0 bz bw]. unfold zvec4_max. simpl.
  apply zvec4_eq; apply Z.max_comm.
Qed.

Theorem zvec4_min_self : forall a : ZVec4,
  zvec4_min a a = a.
Proof.
  intros [ax ay az aw]. unfold zvec4_min. simpl.
  apply zvec4_eq; apply Z.min_id.
Qed.

Theorem zvec4_max_self : forall a : ZVec4,
  zvec4_max a a = a.
Proof.
  intros [ax ay az aw]. unfold zvec4_max. simpl.
  apply zvec4_eq; apply Z.max_id.
Qed.

(** ** Abs Properties *)

Theorem zvec4_abs_nonneg : forall v : ZVec4,
  0 <= zvec4_x (zvec4_abs v) /\ 0 <= zvec4_y (zvec4_abs v) /\
  0 <= zvec4_z (zvec4_abs v) /\ 0 <= zvec4_w (zvec4_abs v).
Proof.
  intros [vx vy vz vw]. unfold zvec4_abs. simpl.
  repeat split; apply Z.abs_nonneg.
Qed.

Theorem zvec4_abs_neg : forall v : ZVec4,
  zvec4_abs (zvec4_neg v) = zvec4_abs v.
Proof.
  intros [vx vy vz vw]. unfold zvec4_abs, zvec4_neg. simpl.
  apply zvec4_eq; apply Z.abs_opp.
Qed.

Theorem zvec4_abs_idempotent : forall v : ZVec4,
  zvec4_abs (zvec4_abs v) = zvec4_abs v.
Proof.
  intros [vx vy vz vw]. unfold zvec4_abs. simpl.
  apply zvec4_eq; apply Z.abs_eq; apply Z.abs_nonneg.
Qed.

(** ** Distance Properties *)

Theorem zvec4_distance_squared_self : forall a : ZVec4,
  zvec4_distance_squared a a = 0.
Proof.
  intros [ax ay az aw].
  unfold zvec4_distance_squared, zvec4_length_squared, zvec4_sub, zvec4_dot.
  simpl. ring.
Qed.

Theorem zvec4_distance_squared_symmetric : forall a b : ZVec4,
  zvec4_distance_squared a b = zvec4_distance_squared b a.
Proof.
  intros [ax ay az aw] [bx by0 bz bw].
  unfold zvec4_distance_squared, zvec4_length_squared, zvec4_sub, zvec4_dot.
  simpl. ring.
Qed.

Theorem zvec4_distance_squared_nonneg : forall a b : ZVec4,
  0 <= zvec4_distance_squared a b.
Proof.
  intros [ax ay az aw] [bx by0 bz bw].
  unfold zvec4_distance_squared, zvec4_length_squared, zvec4_sub, zvec4_dot.
  simpl.
  apply Z.add_nonneg_nonneg; [apply Z.add_nonneg_nonneg; [apply Z.add_nonneg_nonneg |] |]; apply Z.square_nonneg.
Qed.

(** ** Element Sum/Product Properties *)

Theorem zvec4_element_sum_zero :
  zvec4_element_sum zvec4_zero = 0.
Proof.
  unfold zvec4_element_sum, zvec4_zero. simpl. reflexivity.
Qed.

(** * Computational Tests *)

Example zvec4_test_add :
  zvec4_add (mkZVec4 1 2 3 4) (mkZVec4 5 6 7 8) = mkZVec4 6 8 10 12.
Proof. reflexivity. Qed.

Example zvec4_test_dot :
  zvec4_dot (mkZVec4 1 2 3 4) (mkZVec4 5 6 7 8) = 70.
Proof. reflexivity. Qed.

Example zvec4_test_scale :
  zvec4_scale 3 (mkZVec4 2 5 7 11) = mkZVec4 6 15 21 33.
Proof. reflexivity. Qed.

Example zvec4_test_length_sq :
  zvec4_length_squared (mkZVec4 1 2 2 4) = 25.
Proof. reflexivity. Qed.

(** * Notation *)

Notation "a +z4 b" := (zvec4_add a b) (at level 50, left associativity).
Notation "a -z4 b" := (zvec4_sub a b) (at level 50, left associativity).
Notation "s *z4 v" := (zvec4_scale s v) (at level 40, left associativity).
Notation "a .*z4 b" := (zvec4_mul a b) (at level 40, left associativity).
Notation "a ·z4 b" := (zvec4_dot a b) (at level 40, no associativity).
