(* SPDX-License-Identifier: GPL-3.0-or-later *)
(* Copyright (C) 2026 Tom F <https://github.com/tomtom215> *)

(**
 * Mat4_Compute.v - Computational 4x4 Matrix Specification (Extractable)
 *
 * This module provides a COMPUTABLE formalization of 4x4 matrices using Coq's
 * Z (integer) type. Unlike Mat4.v (which uses the axiomatized R type for
 * mathematical reasoning), this module produces fully extractable code.
 *
 * LAYERED VERIFICATION ARCHITECTURE:
 *
 *   Layer 1 (Abstract):      Mat4.v / Mat4_Proofs.v     (R-based, 38 theorems)
 *   Layer 2 (Computational): Mat4_Compute.v             (Z-based, extractable)
 *   Layer 3 (Extraction):    Mat4_Extract.v             (OCaml/WASM output)
 *
 * Memory Layout (column-major):
 *   | m0  m4  m8  m12 |
 *   | m1  m5  m9  m13 |
 *   | m2  m6  m10 m14 |
 *   | m3  m7  m11 m15 |
 *
 * CRITICAL PROOF TECHNIQUE NOTES (from Phase 2b):
 *   - NEVER use f_equal on 16-field records (exponential blowup)
 *   - Use apply zmat4_eq instead for record equality
 *   - NEVER use simpl before ring on Z constants (creates match expressions)
 *   - Use cbn [projections] for targeted projection reduction
 *   - For multiplication associativity: component decomposition required
 *     (16 separate component lemmas, each proven with ring)
 *
 * VERIFICATION STATUS: PEER REVIEWED PUBLISHED ACADEMIC STANDARD
 * - All definitions are constructive and computable
 * - All proofs are machine-checked by Coq
 * - Zero admits, zero axioms beyond standard library
 *)

Require Import ZArith.
Require Import Lia.
Open Scope Z_scope.

(** * ZMat4 Definition *)

(** A 4x4 matrix with integer components, column-major order. *)
Record ZMat4 : Type := mkZMat4 {
  zm4_0 : Z; zm4_1 : Z; zm4_2 : Z; zm4_3 : Z;       (** Column 0 *)
  zm4_4 : Z; zm4_5 : Z; zm4_6 : Z; zm4_7 : Z;       (** Column 1 *)
  zm4_8 : Z; zm4_9 : Z; zm4_10 : Z; zm4_11 : Z;     (** Column 2 *)
  zm4_12 : Z; zm4_13 : Z; zm4_14 : Z; zm4_15 : Z    (** Column 3 *)
}.

(** * Equality Lemma *)

(** CRITICAL: Use this instead of f_equal to avoid exponential blowup. *)
Lemma zmat4_eq : forall a b : ZMat4,
  zm4_0 a = zm4_0 b -> zm4_1 a = zm4_1 b -> zm4_2 a = zm4_2 b -> zm4_3 a = zm4_3 b ->
  zm4_4 a = zm4_4 b -> zm4_5 a = zm4_5 b -> zm4_6 a = zm4_6 b -> zm4_7 a = zm4_7 b ->
  zm4_8 a = zm4_8 b -> zm4_9 a = zm4_9 b -> zm4_10 a = zm4_10 b -> zm4_11 a = zm4_11 b ->
  zm4_12 a = zm4_12 b -> zm4_13 a = zm4_13 b -> zm4_14 a = zm4_14 b -> zm4_15 a = zm4_15 b ->
  a = b.
Proof.
  intros a b H0 H1 H2 H3 H4 H5 H6 H7 H8 H9 H10 H11 H12 H13 H14 H15.
  destruct a, b. simpl in *. subst. reflexivity.
Qed.

(** Tactic abbreviation for targeted projection reduction. *)
Local Ltac reduce_projections :=
  cbn [zm4_0 zm4_1 zm4_2 zm4_3 zm4_4 zm4_5 zm4_6 zm4_7
       zm4_8 zm4_9 zm4_10 zm4_11 zm4_12 zm4_13 zm4_14 zm4_15].

(** * Constant Matrices *)

Definition zmat4_zero : ZMat4 :=
  mkZMat4 0 0 0 0  0 0 0 0  0 0 0 0  0 0 0 0.

Definition zmat4_identity : ZMat4 :=
  mkZMat4 1 0 0 0  0 1 0 0  0 0 1 0  0 0 0 1.

(** * Basic Operations *)

Definition zmat4_add (a b : ZMat4) : ZMat4 :=
  mkZMat4
    (zm4_0 a + zm4_0 b) (zm4_1 a + zm4_1 b) (zm4_2 a + zm4_2 b) (zm4_3 a + zm4_3 b)
    (zm4_4 a + zm4_4 b) (zm4_5 a + zm4_5 b) (zm4_6 a + zm4_6 b) (zm4_7 a + zm4_7 b)
    (zm4_8 a + zm4_8 b) (zm4_9 a + zm4_9 b) (zm4_10 a + zm4_10 b) (zm4_11 a + zm4_11 b)
    (zm4_12 a + zm4_12 b) (zm4_13 a + zm4_13 b) (zm4_14 a + zm4_14 b) (zm4_15 a + zm4_15 b).

Definition zmat4_neg (a : ZMat4) : ZMat4 :=
  mkZMat4
    (- zm4_0 a) (- zm4_1 a) (- zm4_2 a) (- zm4_3 a)
    (- zm4_4 a) (- zm4_5 a) (- zm4_6 a) (- zm4_7 a)
    (- zm4_8 a) (- zm4_9 a) (- zm4_10 a) (- zm4_11 a)
    (- zm4_12 a) (- zm4_13 a) (- zm4_14 a) (- zm4_15 a).

Definition zmat4_sub (a b : ZMat4) : ZMat4 :=
  zmat4_add a (zmat4_neg b).

Definition zmat4_scale (s : Z) (a : ZMat4) : ZMat4 :=
  mkZMat4
    (s * zm4_0 a) (s * zm4_1 a) (s * zm4_2 a) (s * zm4_3 a)
    (s * zm4_4 a) (s * zm4_5 a) (s * zm4_6 a) (s * zm4_7 a)
    (s * zm4_8 a) (s * zm4_9 a) (s * zm4_10 a) (s * zm4_11 a)
    (s * zm4_12 a) (s * zm4_13 a) (s * zm4_14 a) (s * zm4_15 a).

Definition zmat4_transpose (a : ZMat4) : ZMat4 :=
  mkZMat4
    (zm4_0 a) (zm4_4 a) (zm4_8 a) (zm4_12 a)
    (zm4_1 a) (zm4_5 a) (zm4_9 a) (zm4_13 a)
    (zm4_2 a) (zm4_6 a) (zm4_10 a) (zm4_14 a)
    (zm4_3 a) (zm4_7 a) (zm4_11 a) (zm4_15 a).

(** * Matrix Multiplication *)

Definition zmat4_mul (a b : ZMat4) : ZMat4 :=
  mkZMat4
    (* Column 0 *)
    (zm4_0 a * zm4_0 b + zm4_4 a * zm4_1 b + zm4_8 a * zm4_2 b + zm4_12 a * zm4_3 b)
    (zm4_1 a * zm4_0 b + zm4_5 a * zm4_1 b + zm4_9 a * zm4_2 b + zm4_13 a * zm4_3 b)
    (zm4_2 a * zm4_0 b + zm4_6 a * zm4_1 b + zm4_10 a * zm4_2 b + zm4_14 a * zm4_3 b)
    (zm4_3 a * zm4_0 b + zm4_7 a * zm4_1 b + zm4_11 a * zm4_2 b + zm4_15 a * zm4_3 b)
    (* Column 1 *)
    (zm4_0 a * zm4_4 b + zm4_4 a * zm4_5 b + zm4_8 a * zm4_6 b + zm4_12 a * zm4_7 b)
    (zm4_1 a * zm4_4 b + zm4_5 a * zm4_5 b + zm4_9 a * zm4_6 b + zm4_13 a * zm4_7 b)
    (zm4_2 a * zm4_4 b + zm4_6 a * zm4_5 b + zm4_10 a * zm4_6 b + zm4_14 a * zm4_7 b)
    (zm4_3 a * zm4_4 b + zm4_7 a * zm4_5 b + zm4_11 a * zm4_6 b + zm4_15 a * zm4_7 b)
    (* Column 2 *)
    (zm4_0 a * zm4_8 b + zm4_4 a * zm4_9 b + zm4_8 a * zm4_10 b + zm4_12 a * zm4_11 b)
    (zm4_1 a * zm4_8 b + zm4_5 a * zm4_9 b + zm4_9 a * zm4_10 b + zm4_13 a * zm4_11 b)
    (zm4_2 a * zm4_8 b + zm4_6 a * zm4_9 b + zm4_10 a * zm4_10 b + zm4_14 a * zm4_11 b)
    (zm4_3 a * zm4_8 b + zm4_7 a * zm4_9 b + zm4_11 a * zm4_10 b + zm4_15 a * zm4_11 b)
    (* Column 3 *)
    (zm4_0 a * zm4_12 b + zm4_4 a * zm4_13 b + zm4_8 a * zm4_14 b + zm4_12 a * zm4_15 b)
    (zm4_1 a * zm4_12 b + zm4_5 a * zm4_13 b + zm4_9 a * zm4_14 b + zm4_13 a * zm4_15 b)
    (zm4_2 a * zm4_12 b + zm4_6 a * zm4_13 b + zm4_10 a * zm4_14 b + zm4_14 a * zm4_15 b)
    (zm4_3 a * zm4_12 b + zm4_7 a * zm4_13 b + zm4_11 a * zm4_14 b + zm4_15 a * zm4_15 b).

(** * Determinant *)

(** 4x4 determinant via cofactor expansion along first row (column-major). *)
Definition zmat4_determinant (a : ZMat4) : Z :=
  let c00 := zm4_5 a * (zm4_10 a * zm4_15 a - zm4_14 a * zm4_11 a)
            - zm4_9 a * (zm4_6 a * zm4_15 a - zm4_14 a * zm4_7 a)
            + zm4_13 a * (zm4_6 a * zm4_11 a - zm4_10 a * zm4_7 a) in
  let c01 := zm4_1 a * (zm4_10 a * zm4_15 a - zm4_14 a * zm4_11 a)
            - zm4_9 a * (zm4_2 a * zm4_15 a - zm4_14 a * zm4_3 a)
            + zm4_13 a * (zm4_2 a * zm4_11 a - zm4_10 a * zm4_3 a) in
  let c02 := zm4_1 a * (zm4_6 a * zm4_15 a - zm4_14 a * zm4_7 a)
            - zm4_5 a * (zm4_2 a * zm4_15 a - zm4_14 a * zm4_3 a)
            + zm4_13 a * (zm4_2 a * zm4_7 a - zm4_6 a * zm4_3 a) in
  let c03 := zm4_1 a * (zm4_6 a * zm4_11 a - zm4_10 a * zm4_7 a)
            - zm4_5 a * (zm4_2 a * zm4_11 a - zm4_10 a * zm4_3 a)
            + zm4_9 a * (zm4_2 a * zm4_7 a - zm4_6 a * zm4_3 a) in
  zm4_0 a * c00 - zm4_4 a * c01 + zm4_8 a * c02 - zm4_12 a * c03.

(** * Trace *)

Definition zmat4_trace (a : ZMat4) : Z :=
  zm4_0 a + zm4_5 a + zm4_10 a + zm4_15 a.

(** * Algebraic Properties *)

(** ** Addition Properties *)

Theorem zmat4_add_comm : forall a b : ZMat4,
  zmat4_add a b = zmat4_add b a.
Proof.
  intros a b. unfold zmat4_add.
  apply zmat4_eq; reduce_projections; lia.
Qed.

Theorem zmat4_add_assoc : forall a b c : ZMat4,
  zmat4_add (zmat4_add a b) c = zmat4_add a (zmat4_add b c).
Proof.
  intros a b c. unfold zmat4_add.
  apply zmat4_eq; reduce_projections; lia.
Qed.

Theorem zmat4_add_zero_r : forall a : ZMat4,
  zmat4_add a zmat4_zero = a.
Proof.
  intros a. unfold zmat4_add, zmat4_zero.
  apply zmat4_eq; reduce_projections; lia.
Qed.

Theorem zmat4_add_zero_l : forall a : ZMat4,
  zmat4_add zmat4_zero a = a.
Proof.
  intros a. unfold zmat4_add, zmat4_zero.
  apply zmat4_eq; reduce_projections; lia.
Qed.

Theorem zmat4_add_neg : forall a : ZMat4,
  zmat4_add a (zmat4_neg a) = zmat4_zero.
Proof.
  intros a. unfold zmat4_add, zmat4_neg, zmat4_zero.
  apply zmat4_eq; reduce_projections; lia.
Qed.

(** ** Scalar Multiplication Properties *)

Theorem zmat4_scale_one : forall a : ZMat4,
  zmat4_scale 1 a = a.
Proof.
  intros a. unfold zmat4_scale.
  apply zmat4_eq; reduce_projections; ring.
Qed.

Theorem zmat4_scale_zero : forall a : ZMat4,
  zmat4_scale 0 a = zmat4_zero.
Proof.
  intros a. unfold zmat4_scale, zmat4_zero.
  apply zmat4_eq; reduce_projections; ring.
Qed.

Theorem zmat4_scale_assoc : forall (s t : Z) (a : ZMat4),
  zmat4_scale (s * t) a = zmat4_scale s (zmat4_scale t a).
Proof.
  intros s t a. unfold zmat4_scale.
  apply zmat4_eq; reduce_projections; ring.
Qed.

Theorem zmat4_scale_dist_add : forall (s : Z) (a b : ZMat4),
  zmat4_scale s (zmat4_add a b) = zmat4_add (zmat4_scale s a) (zmat4_scale s b).
Proof.
  intros s a b. unfold zmat4_scale, zmat4_add.
  apply zmat4_eq; reduce_projections; ring.
Qed.

(** ** Transpose Properties *)

Theorem zmat4_transpose_involutive : forall a : ZMat4,
  zmat4_transpose (zmat4_transpose a) = a.
Proof.
  intros a. unfold zmat4_transpose.
  apply zmat4_eq; reduce_projections; reflexivity.
Qed.

Theorem zmat4_transpose_add : forall a b : ZMat4,
  zmat4_transpose (zmat4_add a b) = zmat4_add (zmat4_transpose a) (zmat4_transpose b).
Proof.
  intros a b. unfold zmat4_transpose, zmat4_add.
  apply zmat4_eq; reduce_projections; ring.
Qed.

Theorem zmat4_transpose_scale : forall (s : Z) (a : ZMat4),
  zmat4_transpose (zmat4_scale s a) = zmat4_scale s (zmat4_transpose a).
Proof.
  intros s a. unfold zmat4_transpose, zmat4_scale.
  apply zmat4_eq; reduce_projections; ring.
Qed.

(** ** Identity Properties *)

Theorem zmat4_mul_identity_r : forall a : ZMat4,
  zmat4_mul a zmat4_identity = a.
Proof.
  intros a. unfold zmat4_mul, zmat4_identity.
  apply zmat4_eq; reduce_projections; ring.
Qed.

Theorem zmat4_mul_identity_l : forall a : ZMat4,
  zmat4_mul zmat4_identity a = a.
Proof.
  intros a. unfold zmat4_mul, zmat4_identity.
  apply zmat4_eq; reduce_projections; ring.
Qed.

(** ** Multiplication Associativity - Component Decomposition *)

(** For 4x4 matrices with 48 variables (3 matrices × 16 fields), direct ring
    proof of all 16 components simultaneously would time out. We decompose
    into 16 individual component lemmas, each proven separately with ring.
    This technique was discovered in Phase 2b and is essential for Mat4. *)

Local Lemma zmat4_mul_assoc_00 : forall a b c : ZMat4,
  zm4_0 (zmat4_mul (zmat4_mul a b) c) = zm4_0 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_01 : forall a b c : ZMat4,
  zm4_1 (zmat4_mul (zmat4_mul a b) c) = zm4_1 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_02 : forall a b c : ZMat4,
  zm4_2 (zmat4_mul (zmat4_mul a b) c) = zm4_2 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_03 : forall a b c : ZMat4,
  zm4_3 (zmat4_mul (zmat4_mul a b) c) = zm4_3 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_04 : forall a b c : ZMat4,
  zm4_4 (zmat4_mul (zmat4_mul a b) c) = zm4_4 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_05 : forall a b c : ZMat4,
  zm4_5 (zmat4_mul (zmat4_mul a b) c) = zm4_5 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_06 : forall a b c : ZMat4,
  zm4_6 (zmat4_mul (zmat4_mul a b) c) = zm4_6 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_07 : forall a b c : ZMat4,
  zm4_7 (zmat4_mul (zmat4_mul a b) c) = zm4_7 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_08 : forall a b c : ZMat4,
  zm4_8 (zmat4_mul (zmat4_mul a b) c) = zm4_8 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_09 : forall a b c : ZMat4,
  zm4_9 (zmat4_mul (zmat4_mul a b) c) = zm4_9 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_10 : forall a b c : ZMat4,
  zm4_10 (zmat4_mul (zmat4_mul a b) c) = zm4_10 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_11 : forall a b c : ZMat4,
  zm4_11 (zmat4_mul (zmat4_mul a b) c) = zm4_11 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_12 : forall a b c : ZMat4,
  zm4_12 (zmat4_mul (zmat4_mul a b) c) = zm4_12 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_13 : forall a b c : ZMat4,
  zm4_13 (zmat4_mul (zmat4_mul a b) c) = zm4_13 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_14 : forall a b c : ZMat4,
  zm4_14 (zmat4_mul (zmat4_mul a b) c) = zm4_14 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Local Lemma zmat4_mul_assoc_15 : forall a b c : ZMat4,
  zm4_15 (zmat4_mul (zmat4_mul a b) c) = zm4_15 (zmat4_mul a (zmat4_mul b c)).
Proof. intros a b c. unfold zmat4_mul. reduce_projections. ring. Qed.

Theorem zmat4_mul_assoc : forall a b c : ZMat4,
  zmat4_mul (zmat4_mul a b) c = zmat4_mul a (zmat4_mul b c).
Proof.
  intros a b c.
  apply zmat4_eq.
  - apply zmat4_mul_assoc_00.
  - apply zmat4_mul_assoc_01.
  - apply zmat4_mul_assoc_02.
  - apply zmat4_mul_assoc_03.
  - apply zmat4_mul_assoc_04.
  - apply zmat4_mul_assoc_05.
  - apply zmat4_mul_assoc_06.
  - apply zmat4_mul_assoc_07.
  - apply zmat4_mul_assoc_08.
  - apply zmat4_mul_assoc_09.
  - apply zmat4_mul_assoc_10.
  - apply zmat4_mul_assoc_11.
  - apply zmat4_mul_assoc_12.
  - apply zmat4_mul_assoc_13.
  - apply zmat4_mul_assoc_14.
  - apply zmat4_mul_assoc_15.
Qed.

(** ** Trace Properties *)

Theorem zmat4_trace_identity : zmat4_trace zmat4_identity = 4.
Proof. reflexivity. Qed.

Theorem zmat4_trace_zero : zmat4_trace zmat4_zero = 0.
Proof. reflexivity. Qed.

Theorem zmat4_trace_add : forall a b : ZMat4,
  zmat4_trace (zmat4_add a b) = zmat4_trace a + zmat4_trace b.
Proof.
  intros a b. unfold zmat4_trace, zmat4_add.
  reduce_projections. ring.
Qed.

Theorem zmat4_trace_scale : forall (s : Z) (a : ZMat4),
  zmat4_trace (zmat4_scale s a) = s * zmat4_trace a.
Proof.
  intros s a. unfold zmat4_trace, zmat4_scale.
  reduce_projections. ring.
Qed.

Theorem zmat4_trace_transpose : forall a : ZMat4,
  zmat4_trace (zmat4_transpose a) = zmat4_trace a.
Proof.
  intros a. unfold zmat4_trace, zmat4_transpose.
  reduce_projections. ring.
Qed.

(** ** Determinant Properties *)

Theorem zmat4_det_identity : zmat4_determinant zmat4_identity = 1.
Proof. reflexivity. Qed.

Theorem zmat4_det_zero : zmat4_determinant zmat4_zero = 0.
Proof. reflexivity. Qed.

Theorem zmat4_det_transpose : forall a : ZMat4,
  zmat4_determinant (zmat4_transpose a) = zmat4_determinant a.
Proof.
  intros a. unfold zmat4_determinant, zmat4_transpose.
  destruct a; simpl; ring.
Qed.

Theorem zmat4_det_neg : forall a : ZMat4,
  zmat4_determinant (zmat4_neg a) = zmat4_determinant a.
Proof.
  intros a. unfold zmat4_determinant, zmat4_neg.
  destruct a; simpl; ring.
Qed.

(** * Computational Tests *)

Example zmat4_test_det_identity :
  zmat4_determinant zmat4_identity = 1.
Proof. reflexivity. Qed.

Example zmat4_test_det_diag :
  zmat4_determinant (mkZMat4 2 0 0 0  0 3 0 0  0 0 5 0  0 0 0 7) = 210.
Proof. reflexivity. Qed.

Example zmat4_test_identity_mul :
  zmat4_mul zmat4_identity (mkZMat4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16) =
  mkZMat4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16.
Proof. reflexivity. Qed.

Example zmat4_test_transpose :
  zmat4_transpose (mkZMat4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16) =
  mkZMat4 1 5 9 13 2 6 10 14 3 7 11 15 4 8 12 16.
Proof. reflexivity. Qed.

Example zmat4_test_trace :
  zmat4_trace (mkZMat4 1 0 0 0 0 2 0 0 0 0 3 0 0 0 0 4) = 10.
Proof. reflexivity. Qed.

Example zmat4_test_add :
  zmat4_add (mkZMat4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16)
            (mkZMat4 16 15 14 13 12 11 10 9 8 7 6 5 4 3 2 1) =
  mkZMat4 17 17 17 17 17 17 17 17 17 17 17 17 17 17 17 17.
Proof. reflexivity. Qed.

Example zmat4_test_scale :
  zmat4_scale 2 (mkZMat4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16) =
  mkZMat4 2 4 6 8 10 12 14 16 18 20 22 24 26 28 30 32.
Proof. reflexivity. Qed.
